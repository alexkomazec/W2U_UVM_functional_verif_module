//------------------------------------------------------------------------------
// Copyright (c) 2019 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : wb2uart_virtual_sequence_lib.sv
// Developer  : Aleksandar Komazec
// Date       :
// Description:
// Notes      :
//
//------------------------------------------------------------------------------

`ifndef WB2UART_VIRTUAL_SEQUENCE_LIB_SV
`define WB2UART_VIRTUAL_SEQUENCE_LIB_SV

`include "wb2uart_virtual_sequence_base.sv"
`include "wb2uart_virtual_seq_register_access.sv"
`include "wb2uart_virtual_seq_dut_config.sv"
`include "wb2uart_virtual_seq_interrupt_trigger.sv"
`include "wb2uart_virtual_seq_fifo_wr_rd.sv"

`endif // WB2UART_VIRTUAL_SEQUENCE_LIB_SV


