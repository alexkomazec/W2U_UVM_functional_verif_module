//------------------------------------------------------------------------------
// Copyright (c) 2019 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : uart_uvc_tx_seq_lib.sv
// Developer  : Aleksandar Komazec
// Date       :
// Description:
// Notes      :
//
//------------------------------------------------------------------------------

`ifndef UART_UVC_TX_SEQ_LIB_SV
`define UART_UVC_TX_SEQ_LIB_SV

`include "uart_uvc_tx_seq.sv"

`endif // UART_UVC_TX_SEQ_LIB_SV
