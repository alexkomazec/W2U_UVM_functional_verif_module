//------------------------------------------------------------------------------
// Copyright (c) 2019 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : wb2uart_common.sv
// Developer  : Aleksandar Komazec
// Date       :
// Description: 
// Notes      : 
//
//------------------------------------------------------------------------------

`ifndef WB2UART_COMMON_SV
`define WB2UART_COMMON_SV

int virtual_Sequence_register_access_time_out = 99999999;


`endif // WB2UART_COMMON_SV
